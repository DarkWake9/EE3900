
V1 in 0 SIN (0 12 5k 0 0)
R0 in 1 1
C1 1 0 1.64m ic=0
L2 1 2 4.29m
C3 2 0 5.31m ic=0
L4 2 3 4.29m
C5 X 0 1.64m ic=0
RL X 0 1
V2 out

.control
tran 1e-9 10u uic
plot  v(X)
wrdata e5.3b.txt v(X)
.endc

.end
