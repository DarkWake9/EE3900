* Output After Switching

R1  X    0    1

C1  X    0    1u    ic=0

R2  X    1    2

V2  1    0    dc	2V


.control
tran    100n    10u    uic

run
wrdata    e4.txt    v(X)
set color0 = white
set color1 = black
plot  v(X)
hardcopy ../figs/e4.7.pdf v(X)
.endc

.end
